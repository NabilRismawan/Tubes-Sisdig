library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


ENTITY LUTArcCos IS
    PORT (
        masukan : IN STD_LOGIC_VECTOR (31 downto 0); -- Input: 32 bit
        keluaran : OUT STD_LOGIC_VECTOR (15 downto 0) -- Output: 16 bite
			);
END LUTArcCos;

ARCHITECTURE Behavioral OF LUTArcCos IS 
BEGIN 
    Process (masukan) is
    BEGIN 
        -- keluaran <= (others => "0");
        case masukan is
            -- input 32bit ke biner 16 bit
            when "11111111100000000000000000000000" => keluaran <= "1011010000000000"; -- input = -1, output = 180 derajat
            when "11111111011111001111010111010011" => keluaran <= "1010101111100010"; -- -0.99
            when "11111111011110010011011010011010" => keluaran <= "1010100000100010"; -- -0.98 
            when "11111111011101111010101100101000" => keluaran <= "1010011111101100"; -- -0.97
            when "11111111011100111010100011001100" => keluaran <= "1010011100111100"; -- -0.96
            when "11111111011011111110101001010001" => keluaran <= "1010011011010111"; -- -0.95
            when "11111111011011000110111111100001" => keluaran <= "1010011001000101"; -- -0.94
            when "11111111011010001111001110001000" => keluaran <= "1010010111100000"; -- -0.93
            when "11111111011001010110101111110101" => keluaran <= "1010010101110110"; -- -0.92
            when "11111111011000011110100011100000" => keluaran <= "1010010011110000"; -- -0.91
            when "11111111010111100110011011010100" => keluaran <= "1010010010100000"; -- -0.9
            when "11111111010110101110010011010010" => keluaran <= "1010010001011101"; -- -0.89
            when "11111111010101110110000011111010" => keluaran <= "1010010000101101"; -- -0.88	
            when "11111111010101000001011110101000" => keluaran <= "1010001111111101"; -- -0.87
            when "11111111010011101010110111011011" => keluaran <= "1010001111010001"; -- -0.86	
            when "11111111010010110110110111001001" => keluaran <= "1010001110001100"; -- -0.85	
            when "11111111010010000010001010110011" => keluaran <= "1010001101011011"; -- -0.84
            when "11111111010001001101111110011111" => keluaran <= "1010001100100001"; -- -0.83	
            when "11111111010000011001110110011011" => keluaran <= "1010001011111010"; -- -0.82	
            when "11111111001111100101101010111111" => keluaran <= "1010001011011101"; -- -0.81
            when "11111111001110110001011110110100" => keluaran <= "1010001010110101"; -- -0.8	
            when "11111111001101111101000011011010" => keluaran <= "1010001010011011"; -- -0.79
            when "11111111001101001000100110111000" => keluaran <= "1010001001111100"; -- -0.78	
            when "11111111001100010100001101100000" => keluaran <= "1010001001100001"; -- -0.77	
            when "11111111001011100000001010000001" => keluaran <= "1010001001001000"; -- -0.76
            when "11111111001010101100000011011110" => keluaran <= "1010001000110010"; -- -0.75
            when "11111111001001111000000110001110" => keluaran <= "1010001000011000"; -- -0.74
            when "11111111001001000100001100000000" => keluaran <= "1010000111111101"; -- -0.73	
            when "11111111001000010000010010011110" => keluaran <= "1010000111101001"; -- -0.72
            when "11111111000111011100100010000010" => keluaran <= "1010000111010101"; -- -0.71
            when "11111111000110101000110001000000" => keluaran <= "1010000110111111"; -- -0.70
            when "11111111000101110101000010111010" => keluaran <= "1010000110101101"; -- -0.69
            when "11111111000101000001010110100001" => keluaran <= "1010000110011001"; -- -0.68
            when "11111111000011001101110110010000" => keluaran <= "1010000110000111"; -- -0.67
            when "11111111000010011010100001001100" => keluaran <= "1010000101110100"; -- -0.66
            when "11111111000001100111011101001001" => keluaran <= "1010000101100001"; -- -0.65
            when "11111111000000110011110101011110" => keluaran <= "1010000101001000"; -- -0.64
            when "11111110111111111100100100010100" => keluaran <= "1010000100110100"; -- -0.63
            when "11111110111111010001010000000001" => keluaran <= "1010000100011000"; -- -0.62
            when "11111110111110011101101011010110" => keluaran <= "1010000011111101"; -- -0.61
            when "11111110111101101010011011101101" => keluaran <= "1010000011101000"; -- -0.60
            when "11111110111100110111000100001001" => keluaran <= "1010000011010010"; -- -0.59
            when "11111110111011111111101010011111" => keluaran <= "1010000010111111"; -- -0.58
            when "11111110111011001000011010100011" => keluaran <= "1010000010101101"; -- -0.57
            when "11111110111010010001000000010001" => keluaran <= "1010000010011000"; -- -0.56
            when "11111110111001100001101101001010" => keluaran <= "1010000010000110"; -- -0.55
            when "11111110111000101010010111110010" => keluaran <= "1010000001110101"; -- -0.54
            when "11111110110111110011001010111000" => keluaran <= "1010000001100101"; -- -0.53
            when "11111110110111000000000000010111" => keluaran <= "1010000001010101"; -- -0.52
            when "11111110110110001001010110011100" => keluaran <= "1010000001000100"; -- -0.51
            when "11111110110101010010101010111001" => keluaran <= "1010000000110000"; -- -0.50
            when "11111110110100011100011011110101" => keluaran <= "1010000000011101"; -- -0.49
            when "11111110110011100110011110101011" => keluaran <= "1010000000001001"; -- -0.48
            when "11111110110010110000110111010001" => keluaran <= "1001111111110000"; -- -0.47
            when "11111110110001111111010011001010" => keluaran <= "1001111111100011"; -- -0.46
            when "11111110110001001001101110011011" => keluaran <= "1001111111010110"; -- -0.45
            when "11111110110000010011110011101100" => keluaran <= "1001111111001001"; -- -0.44
            when "11111110101111011101111110100000" => keluaran <= "1001111110111100"; -- -0.43
            when "11111110101110101011110001110001" => keluaran <= "1001111110101111"; -- -0.42
            when "11111110101101110101110110100000" => keluaran <= "1001111110011101"; -- -0.41
            when "11111110101101000000001000011111" => keluaran <= "1001111110001111"; -- -0.40
            when "11111110101100001010011011111110" => keluaran <= "1001111101111101"; -- -0.39
            when "11111110101011010100111111101001" => keluaran <= "1001111101101110"; -- -0.38
            when "11111110101010100011110010011000" => keluaran <= "1001111101011100"; -- -0.37
            when "11111110101001110010101000110111" => keluaran <= "1001111101001101"; -- -0.36
            when "11111110101001000001110101011110" => keluaran <= "1001111100111101"; -- -0.35
            when "11111110101000010001000001101000" => keluaran <= "1001111100101101"; -- -0.34
            when "11111110100111100000000111010101" => keluaran <= "1001111100011101"; -- -0.33
            when "11111110100110110011001100110000" => keluaran <= "1001111100001110"; -- -0.32
            when "11111110100110000010011001100110" => keluaran <= "1001111011111100"; -- -0.31
            when "11111110100101010001110011110001" => keluaran <= "1001111011101100"; -- -0.30
            when "11111110100100100001000111111001" => keluaran <= "1001111011011100"; -- -0.29
            when "11111110100011110000011111100110" => keluaran <= "1001111011001100"; -- -0.28
            when "11111110100011000000000000010000" => keluaran <= "1001111010111100"; -- -0.27
            when "11111110100010010000100110110111" => keluaran <= "1001111010101101"; -- -0.26
            when "11111110100001100001010011000001" => keluaran <= "1001111010011101"; -- -0.25
            when "11111110100000110001101111001000" => keluaran <= "1001111010001110"; -- -0.24
            when "11111110011111111110001000111101" => keluaran <= "1001111001111111"; -- -0.23
            when "11111110011111001110100010010010" => keluaran <= "1001111001101111"; -- -0.22
            when "11111110011110011110111100001011" => keluaran <= "1001111001011111"; -- -0.21
            when "11111110011101101111010010100011" => keluaran <= "1001111001001111"; -- -0.20
            when "11111110011100111111100100110101" => keluaran <= "1001111000111111"; -- -0.19
            when "11111110011011110000000001000011" => keluaran <= "1001111000101111"; -- -0.18
            when "11111110011011000000010110010001" => keluaran <= "1001111000011111"; -- -0.17
            when "11111110011010010000101011010100" => keluaran <= "1001111000001111"; -- -0.16
            when "11111110011001100000111111110110" => keluaran <= "1001110111111111"; -- -0.15
            when "11111110011000110001010100010101" => keluaran <= "1001110111101111"; -- -0.14
            when "11111110010111111101101000010000" => keluaran <= "1001110111011111"; -- -0.13
            when "11111110010111001110000000001010" => keluaran <= "1001110111001111"; -- -0.12
            when "11111110010110011110010011011001" => keluaran <= "1001110110111111"; -- -0.11
            when "11111110010101101110100111001001" => keluaran <= "1001110110101111"; -- -0.10
            when "11111110010100111110111010111101" => keluaran <= "1001110110011111"; -- -0.09
            when "11111110010011101111001110101010" => keluaran <= "1001110110001111"; -- -0.08
            when "11111110010010111110111111011011" => keluaran <= "1001110101111111"; -- -0.07
            when "11111110010010001110110101001000" => keluaran <= "1001110101101111"; -- -0.06
            when "11111110010001011111001011000010" => keluaran <= "1001110101011111"; -- -0.05
            when "11111110010000101111011111110100" => keluaran <= "1001110101001111"; -- -0.04
            when "11111110001111111111110100110001" => keluaran <= "1001110100111111"; -- -0.03
            when "11111110001111001111100011110000" => keluaran <= "1001110100101111"; -- -0.02
            when "11111110001110011111110010100001" => keluaran <= "1001110100011111"; -- -0.01
            when "00000000000000000000000000000000" => keluaran <= "1001110100001111"; --  0.00
            when "00111111011111110000010000011000" => keluaran <= "1001110011111111"; --  0.01
            when "00111111011111100000100000111000" => keluaran <= "1001110011101111"; --  0.02
            when "00111111011111010000110001010000" => keluaran <= "1001110011011111"; --  0.03
            when "00111111011111000001000001101000" => keluaran <= "1001110011001111"; --  0.04
            when "00111111011110110001010010001000" => keluaran <= "1001110010111111"; --  0.05
            when "00111111011110100001100100100000" => keluaran <= "1001110010101111"; --  0.06
            when "00111111011110010001110111100000" => keluaran <= "1001110010011111"; --  0.07
            when "00111111011110000010001001011000" => keluaran <= "1001110010001111"; --  0.08
            when "00111111011101110010011011110000" => keluaran <= "1001110001111111"; --  0.09
            when "00111111011101100010101100101000" => keluaran <= "1001110001101111"; --  0.10
            when "00111111011101010010111101011000" => keluaran <= "1001110001011111"; --  0.11
            when "00111111011101000011001110110000" => keluaran <= "1001110001001111"; --  0.12
            when "00111111011100110011011110001000" => keluaran <= "1001110000111111"; --  0.13
            when "00111111011100100011101111100000" => keluaran <= "1001110000101111"; --  0.14
            when "00111111011011110011111101011000" => keluaran <= "1001110000011111"; --  0.15
            when "00111111011011100011101011110000" => keluaran <= "1001110000001111"; --  0.16
            when "00111111011011010011011010001000" => keluaran <= "1001101111111111"; --  0.17
            when "00111111011011000011001000100000" => keluaran <= "1001101111101111"; --  0.18
            when "00111111011010110010110110111000" => keluaran <= "1001101111011111"; --  0.19
            when "00111111011010100010100101010000" => keluaran <= "1001101111001111"; --  0.20
            when "00111111011010010010010011101000" => keluaran <= "1001101110111111"; --  0.21
            when "00111111011010000010000010000000" => keluaran <= "1001101110101111"; --  0.22
            when "00111111011001110001110000011000" => keluaran <= "1001101110011111"; --  0.23
            when "00111111011001100001100000110000" => keluaran <= "1001101110001111"; --  0.24
            when "00111111011001010001010011001000" => keluaran <= "1001101101111111"; --  0.25
            when "00111111011001000001000100100000" => keluaran <= "1001101101101111"; --  0.26
            when "00111111011000110000110110111000" => keluaran <= "1001101101011111"; --  0.27
            when "00111111011000100000101001010000" => keluaran <= "1001101101001111"; --  0.28
            when "00111111011000010000011111101000" => keluaran <= "1001101100111111"; --  0.29
            when "00111111010111110000010100000000" => keluaran <= "1001101100101111"; --  0.30
            when "00111111010111100000001010011000" => keluaran <= "1001101100011111"; --  0.31
            when "00111111010111010000000000110000" => keluaran <= "1001101100001111"; --  0.32
            when "00111111010111000000010111001000" => keluaran <= "1001101011111111"; --  0.33
            when "00111111010110110000001101111000" => keluaran <= "1001101011101111"; --  0.34
            when "00111111010110100000000011110000" => keluaran <= "1001101011011111"; --  0.35
            when "00111111010110010000011010001000" => keluaran <= "1001101011001111"; --  0.36
            when "00111111010110000000001111111000" => keluaran <= "1001101010111111"; --  0.37
            when "00111111010101110000000101110000" => keluaran <= "1001101010101111"; --  0.38
            when "00111111010101100000011011101000" => keluaran <= "1001101010001111"; --  0.39
            when "00111111010101010000010001110000" => keluaran <= "1001101001111111"; --  0.40
            when "00111111010101000000001011101000" => keluaran <= "1001101001101111"; --  0.41
            when "00111111010100110000000010100000" => keluaran <= "1001101001011111"; --  0.42
            when "00111111010100100000011001011000" => keluaran <= "1001101001001111"; --  0.43
            when "00111111010100010000010000001000" => keluaran <= "1001101000111111"; --  0.44
            when "00111111010011110000000110111000" => keluaran <= "1001101000101111"; --  0.45
            when "00111111010011100000011101110000" => keluaran <= "1001101000011111"; --  0.46
            when "00111111010011010000010100100000" => keluaran <= "1001101000001111"; --  0.47
            when "00111111010011000000001111000000" => keluaran <= "1001100111111111"; --  0.48
            when "00111111010010110000000110010000" => keluaran <= "1001100111101111"; --  0.49
            when "00111111010010100000000001100000" => keluaran <= "1001100111011111"; --  0.50
            when "00111111010010010000011100110000" => keluaran <= "1001100111001111"; --  0.51
            when "00111111010010000000010111011000" => keluaran <= "1001100110111111"; --  0.52
            when "00111111010001110000010010001000" => keluaran <= "1001100110101111"; --  0.53
            when "00111111010001100000001100111000" => keluaran <= "1001100110011111"; --  0.54
            when "00111111010001010000001000001000" => keluaran <= "1001100110001111"; --  0.55
            when "00111111010001000000000011100000" => keluaran <= "1001100101111111"; --  0.56
            when "00111111010000110000000010111000" => keluaran <= "1001100101101111"; --  0.57
            when "00111111010000100000000110010000" => keluaran <= "1001100101011111"; --  0.58
            when "00111111010000010000001001101000" => keluaran <= "1001100101001111"; --  0.59
            when "00111111010000000000001101000000" => keluaran <= "1001100100111111"; --  0.60
            when "00111110111111110000010000011000" => keluaran <= "1001100100101111"; --  0.61
            when "00111110111111100000010000010000" => keluaran <= "1001100100011111"; --  0.62
            when "00111110111111010000010000001000" => keluaran <= "1001100100001111"; --  0.63
            when "00111110111111000000010000000000" => keluaran <= "1001100011111111"; --  0.64
            when "00111110111110110000010000011000" => keluaran <= "1001100011101111"; --  0.65
            when "00111110111110100000010000100000" => keluaran <= "1001100011011111"; --  0.66
            when "00111110111110010000010000101000" => keluaran <= "1001100011001111"; --  0.67
            when "00111110111110000000010000110000" => keluaran <= "1001100010111111"; --  0.68
            when "00111110111101110000010000111000" => keluaran <= "1001100010101111"; --  0.69
            when "00111110111101100000010001000000" => keluaran <= "1001100010011111"; --  0.70
            when "00111110111101010000010001001000" => keluaran <= "1001100010001111"; --  0.71
            when "00111110111101000000010001010000" => keluaran <= "1001100001111111"; --  0.72
            when "00111110111100110000010001011000" => keluaran <= "1001100001101111"; --  0.73
            when "00111110111100100000010001100000" => keluaran <= "1001100001011111"; --  0.74
            when "00111110111100010000010001101000" => keluaran <= "1001100001001111"; --  0.75
            when "00111110111100000000010001110000" => keluaran <= "1001100000111111"; --  0.76
            when "00111110111011110000010001111000" => keluaran <= "1001100000101111"; --  0.77
            when "00111110111011100000010010000000" => keluaran <= "1001100000011111"; --  0.78
            when "00111110111011010000010010001000" => keluaran <= "1001100000001111"; --  0.79
            when "00111110111011000000010010010000" => keluaran <= "1001011111111111"; --  0.80
            when "00111110111010110000010010011000" => keluaran <= "1001011111101111"; --  0.81
            when "00111110111010100000010010100000" => keluaran <= "1001011111011111"; --  0.82
            when "00111110111010010000010010101000" => keluaran <= "1001011111001111"; --  0.83
            when "00111110111010000000010010110000" => keluaran <= "1001011110111111"; --  0.84
            when "00111110111001110000010010111000" => keluaran <= "1001011110101111"; --  0.85
            when "00111110111001100000010011000000" => keluaran <= "1001011110011111"; --  0.86
            when "00111110111001010000010011001000" => keluaran <= "1001011110001111"; --  0.87
            when "00111110111001000000010011010000" => keluaran <= "1001011101111111"; --  0.88
            when "00111110111000110000010011011000" => keluaran <= "1001011101101111"; --  0.89
            when "00111110111000100000010011100000" => keluaran <= "1001011101011111"; --  0.90
            when "00111110111000010000010011101000" => keluaran <= "1001011101001111"; --  0.91
            when "00111110110111110000010100000000" => keluaran <= "1001011100111111"; --  0.92
            when "00111110110111100000010100001000" => keluaran <= "1001011100101111"; --  0.93
            when "00111110110111010000010100010000" => keluaran <= "1001011100011111"; --  0.94
            when "00111110110111000000010100011000" => keluaran <= "1001011100001111"; --  0.95
            when "00111110110110110000010100100000" => keluaran <= "1001011100001111"; --  0.96
            when "00111110110110100000010100101000" => keluaran <= "1001010000101111"; --  0.97
            when "00111110110110010000010100110000" => keluaran <= "1001001101101111"; --  0.98
            when "00111110110110000000010100111000" => keluaran <= "1001001100101111"; --  0.99
            when "00111111100000000000000000000000" => keluaran <= "1001001100001111"; --  1.00
            when others => keluaran <= "0000000000000000";            
        end case;
    end process;
end Behavioral;

-- Arc Cosine	Hasil (in radian)	Hexadecimal	Degree
-- -1	3.141592654	102944	180
-- -0.99	3.00005318	98306	171.8903855
-- -0.98	2.941257811	96379	168.521659
-- -0.97	2.896027136	94897	165.9301323
-- -0.96	2.857798544	93644	163.7397953
-- -0.95	2.824032224	92538	161.8051277
-- -0.94	2.793426632	91535	160.0515564
-- -0.93	2.765209171	90610	158.434815
-- -0.92	2.738876812	89748	156.9260819
-- -0.91	2.714080389	88935	155.5053515
-- -0.9	2.690565842	88164	154.1580672
-- -0.89	2.668141496	87430	152.8732469
-- -0.88	2.646658527	86726	151.6423634
-- -0.87	2.625998647	86049	150.4586395
-- -0.86	2.606065999	85396	149.3165829
-- -0.85	2.586781621	84764	148.2116694
-- -0.84	2.568079549	84151	147.1401196
-- -0.83	2.549904011	83555	146.098738
-- -0.82	2.532207346	82975	145.0847938
-- -0.81	2.514948442	82410	144.0959314
-- -0.8	2.498091545	81857	143.1301024
-- -0.79	2.481605324	81317	142.1855115
-- -0.78	2.465462144	80788	141.2605754
-- -0.77	2.449637478	80270	140.3538889
-- -0.76	2.434109442	79761	139.4641979
-- -0.75	2.418858406	79261	138.5903779
-- -0.74	2.403866685	78770	137.7314156
-- -0.73	2.389118277	78287	136.8863941
-- -0.72	2.374598646	77811	136.0544804
-- -0.71	2.360294536	77342	135.2349153
-- -0.7	2.346193823	76880	134.427004
-- -0.69	2.33228538	76424	133.6301089
-- -0.68	2.318558961	75975	132.843643
-- -0.67	2.305005114	75530	132.0670648
-- -0.66	2.291615088	75092	131.2998728
-- -0.65	2.278380764	74658	130.5416019
-- -0.64	2.265294592	74229	129.7918195
-- -0.63	2.252349538	73805	129.0501225
-- -0.62	2.23953903	73385	128.3161345
-- -0.61	2.226856918	72970	127.589503
-- -0.6	2.214297436	72558	126.8698976
-- -0.59	2.201855168	72150	126.1570082
-- -0.58	2.189525017	71746	125.4505426
-- -0.57	2.177302182	71346	124.7502258
-- -0.56	2.165182127	70949	124.0557977
-- -0.55	2.153160565	70555	123.367013
-- -0.54	2.141233436	70164	122.6836388
-- -0.53	2.129396892	69776	122.0054548
-- -0.52	2.117647277	69391	121.3322515
-- -0.51	2.105981117	69009	120.6638297
-- -0.5	2.094395102	68629	120
-- -0.49	2.08288608	68252	119.3405816
-- -0.48	2.071451039	67877	118.685402
-- -0.47	2.060087105	67505	118.0342965
-- -0.46	2.048791525	67135	117.3871075
-- -0.45	2.037561666	66767	116.743684
-- -0.44	2.026395	66401	116.1038811
-- -0.43	2.015289104	66037	115.4675601
-- -0.42	2.004241647	65675	114.8345875
-- -0.41	1.993250389	65315	114.2048348
-- -0.4	1.982313173	64956	113.5781785
-- -0.39	1.971427919	64600	112.9544994
-- -0.38	1.960592623	64245	112.3336827
-- -0.37	1.949805347	63891	111.7156173
-- -0.36	1.93906422	63539	111.100196
-- -0.35	1.92836743	63189	110.4873151
-- -0.34	1.917713224	62840	109.8768741
-- -0.33	1.907099902	62492	109.2687755
-- -0.32	1.896525814	62145	108.6629249
-- -0.31	1.885989359	61800	108.0592305
-- -0.3	1.875488981	61456	107.4576031
-- -0.29	1.865023165	61113	106.857956
-- -0.28	1.854590436	60771	106.2602047
-- -0.27	1.844189358	60430	105.6642669
-- -0.26	1.83381853	60091	105.0700621
-- -0.25	1.823476582	59752	104.4775122
-- -0.24	1.813162178	59414	103.8865404
-- -0.23	1.80287401	59077	103.2970717
-- -0.22	1.792610797	58740	102.709033
-- -0.21	1.782371287	58405	102.1223522
-- -0.2	1.772154248	58070	101.536959
-- -0.19	1.761958473	57736	100.9527842
-- -0.18	1.751782778	57402	100.3697598
-- -0.17	1.741625996	57070	99.78781906
-- -0.16	1.73148698	56737	99.20689622
-- -0.15	1.7213646	56406	98.62692656
-- -0.14	1.711257742	56074	98.04784625
-- -0.13	1.701165306	55744	97.46959232
-- -0.12	1.691086209	55414	96.89210258
-- -0.11	1.681019377	55084	96.31531557
-- -0.1	1.670963748	54754	95.73917048
-- -0.09	1.660918272	54425	95.16360709
-- -0.08	1.650881907	54096	94.58856574
-- -0.07	1.64085362	53767	94.01398722
-- -0.06	1.630832385	53439	93.43981277
-- -0.05	1.620817184	53111	92.86598398
-- -0.04	1.610807001	52783	92.29244278
-- -0.03	1.600800829	52455	91.71913132
-- -0.02	1.59079766	52127	91.145992
-- -0.01	1.580796493	51800	90.57296734
-- 0	1.570796327	51472	90
-- 0.01	1.56079616	51144	89.42703266
-- 0.02	1.550794993	50816	88.854008
-- 0.03	1.540791825	50489	88.28086868
-- 0.04	1.530785652	50161	87.70755722
-- 0.05	1.52077547	49833	87.13401602
-- 0.06	1.510760268	49505	86.56018723
-- 0.07	1.500739034	49176	85.98601278
-- 0.08	1.490710747	48848	85.41143426
-- 0.09	1.480674382	48519	84.83639291
-- 0.1	1.470628906	48190	84.26082952
-- 0.11	1.460573277	47860	83.68468443
-- 0.12	1.450506444	47530	83.10789742
-- 0.13	1.440427347	47200	82.53040768
-- 0.14	1.430334912	46869	81.95215375
-- 0.15	1.420228054	46538	81.37307344
-- 0.16	1.410105674	46206	80.79310378
-- 0.17	1.399966658	45874	80.21218094
-- 0.18	1.389809876	45541	79.63024019
-- 0.19	1.37963418	45208	79.0472158
-- 0.2	1.369438406	44874	78.46304097
-- 0.21	1.359221367	44539	77.87764776
-- 0.22	1.348981856	44203	77.29096701
-- 0.23	1.338718644	43867	76.70292825
-- 0.24	1.328430476	43530	76.11345964
-- 0.25	1.318116072	43192	75.52248781
-- 0.26	1.307774124	42853	74.92993786
-- 0.27	1.297403295	42513	74.33573315
-- 0.28	1.287002218	42172	73.73979529
-- 0.29	1.276569489	41831	73.14204398
-- 0.3	1.266103673	41488	72.54239688
-- 0.31	1.255603294	41144	71.94076951
-- 0.32	1.24506684	40798	71.33707512
-- 0.33	1.234492752	40452	70.73122451
-- 0.34	1.223879429	40104	70.12312593
-- 0.35	1.213225223	39755	69.51268489
-- 0.36	1.202528433	39404	68.89980398
-- 0.37	1.191787306	39052	68.28438272
-- 0.38	1.18100003	38699	67.66631734
-- 0.39	1.170164734	38344	67.0455006
-- 0.4	1.159279481	37987	66.42182152
-- 0.41	1.148342265	37629	65.7951652
-- 0.42	1.137351007	37269	65.16541251
-- 0.43	1.12630355	36907	64.53243986
-- 0.44	1.115197653	36543	63.89611886
-- 0.45	1.104030988	36177	63.25631605
-- 0.46	1.092801128	35809	62.6128925
-- 0.47	1.081505549	35439	61.96570347
-- 0.48	1.070141614	35066	61.31459799
-- 0.49	1.058706574	34692	60.65941842
-- 0.5	1.047197551	34315	60
-- 0.51	1.035611537	33935	59.33617026
-- 0.52	1.023945376	33553	58.6677485
-- 0.53	1.012195761	33168	57.99454517
-- 0.54	1.000359217	32780	57.31636115
-- 0.55	0.988432089	32389	56.63298703
-- 0.56	0.976410527	31995	55.94420226
-- 0.57	0.964290472	31598	55.24977425
-- 0.58	0.952067636	31197	54.54945736
-- 0.59	0.939737486	30793	53.8429918
-- 0.6	0.927295218	30386	53.13010235
-- 0.61	0.914735736	29974	52.41049704
-- 0.62	0.902053624	29558	51.68386553
-- 0.63	0.889243115	29139	50.94987746
-- 0.64	0.876298061	28715	50.2081805
-- 0.65	0.86321189	28286	49.45839813
-- 0.66	0.849977566	27852	48.70012721
-- 0.67	0.836587539	27413	47.9329352
-- 0.68	0.823033692	26969	47.15635696
-- 0.69	0.809307274	26519	46.36989113
-- 0.7	0.79539883	26064	45.572996
-- 0.71	0.781298117	25602	44.76508467
-- 0.72	0.766994008	25133	43.94551956
-- 0.73	0.752474376	24657	43.11360595
-- 0.74	0.737725968	24174	42.26858443
-- 0.75	0.722734248	23683	41.40962211
-- 0.76	0.707483212	23183	40.53580211
-- 0.77	0.691955175	22674	39.64611115
-- 0.78	0.67613051	22155	38.7394246
-- 0.79	0.659987329	21626	37.81448851
-- 0.8	0.643501109	21086	36.86989765
-- 0.81	0.626644212	20534	35.90406858
-- 0.82	0.609385308	19968	34.91520625
-- 0.83	0.591688642	19388	33.901262
-- 0.84	0.573513104	18793	32.85988038
-- 0.85	0.554811033	18180	31.78833062
-- 0.86	0.535526654	17548	30.68341711
-- 0.87	0.515594006	16895	29.5413605
-- 0.88	0.494934126	16218	28.35763658
-- 0.89	0.473451157	15514	27.12675312
-- 0.9	0.451026812	14779	25.84193276
-- 0.91	0.427512265	14009	24.49464847
-- 0.92	0.402715842	13196	23.07391807
-- 0.93	0.376383482	12333	21.56518502
-- 0.94	0.348166021	11409	19.94844359
-- 0.95	0.317560429	10406	18.19487234
-- 0.96	0.283794109	9299	16.26020471
-- 0.97	0.245565518	8047	14.06986775
-- 0.98	0.200334842	6565	11.47834095
-- 0.99	0.141539473	4638	8.109614456
-- 1	0	0	0
