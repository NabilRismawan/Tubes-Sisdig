-- tes upload github