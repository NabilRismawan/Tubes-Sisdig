-- tes upload github tes tes