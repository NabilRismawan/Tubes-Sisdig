library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


ENTITY LUTArcCos IS
    PORT (
        masukan : IN STD_LOGIC_VECTOR (31 downto 0); -- Input: 32 bit
        keluaran : OUT STD_LOGIC_VECTOR (15 downto 0) -- Output: 16 bit
        -- valid : OUT std_logic -- Signal to indicate if the output is valid
			);
END LUTArcCos;

ARCHITECTURE Behavioral OF LUTArcCos IS 
BEGIN 
    Process (masukan) is
    BEGIN 
        -- keluaran <= (others => "0");
        case masukan is
            -- input 32bit ke biner 16 bit
            when "11111111100000000000000000000000" => keluaran <= "0000000010110100"; -- input = -1, output = 180 derajat
            when "11111111011111001111010111010011" => keluaran <= ""; -- -0.99
            when "11111111011110010011011010011010" => keluaran <= ""; -- -0.98 
            when "11111111011101111010101100101000" => keluaran <= ""; -- -0.97
            when "11111111011100111010100011001100" => keluaran <= ""; -- -0.96
            when "11111111011011111110101001010001" => keluaran <= ""; -- -0.95
            when "11111111011011000110111111100001" => keluaran <= ""; -- -0.94
            when "11111111011010001111001110001000" => keluaran <= ""; -- -0.93
            when "11111111011001010110101111110101" => keluaran <= ""; -- -0.92
            when "11111111011000011110100011100000" => keluaran <= ""; -- -0.91
            when "11111111010111100110011011010100" => keluaran <= ""; -- -0.9
            when "11111111010110101110010011010010" => keluaran <= ""; -- -0.89
            when "11111111010101110110000011111010" => keluaran <= ""; -- -0.88	
            when "11111111010101000001011110101000" => keluaran <= ""; -- -0.87
            when "11111111010011101010110111011011" => keluaran <= ""; -- -0.86	
            when "11111111010010110110110111001001" => keluaran <= ""; -- -0.85	
            when "11111111010010000010001010110011" => keluaran <= ""; -- -0.84
            when "11111111010001001101111110011111" => keluaran <= ""; -- -0.83	
            when "11111111010000011001110110011011" => keluaran <= ""; -- -0.82	
            when "11111111001111100101101010111111" => keluaran <= ""; -- -0.81
            when "11111111001110110001011110110100" => keluaran <= ""; -- -0.8	
            when "11111111001101111101000011011010" => keluaran <= ""; -- -0.79
            when "11111111001101001000100110111000" => keluaran <= ""; -- -0.78	
            when "11111111001100010100001101100000" => keluaran <= ""; -- -0.77	
            when "11111111001011100000001010000001" => keluaran <= ""; -- -0.76
            when "11111111001010101100000011011110" => keluaran <= ""; -- -0.75
            when "11111111001001111000000110001110" => keluaran <= ""; -- -0.74
            when "11111111001001000100001100000000" => keluaran <= ""; -- -0.73	
            when "11111111001000010000010010011110" => keluaran <= ""; -- -0.72
            when "11111111000111011100100010000010" => keluaran <= ""; -- -0.71
            when "11111111000110101000110001000000" => keluaran <= ""; -- -0.70
            when "11111111000101110101000010111010" => keluaran <= ""; -- -0.69
            when "11111111000101000001010110100001" => keluaran <= ""; -- -0.68
            when "11111111000011001101110110010000" => keluaran <= ""; -- -0.67
            when "11111111000010011010100001001100" => keluaran <= ""; -- -0.66
            when "11111111000001100111011101001001" => keluaran <= ""; -- -0.65
            when "11111111000000110011110101011110" => keluaran <= ""; -- -0.64
            when "11111110111111111100100100010100" => keluaran <= ""; -- -0.63
            when "11111110111111010001010000000001" => keluaran <= ""; -- -0.62
            when "11111110111110011101101011010110" => keluaran <= ""; -- -0.61
            when "11111110111101101010011011101101" => keluaran <= ""; -- -0.60
            when "11111110111100110111000100001001" => keluaran <= ""; -- -0.59
            when "11111110111011111111101010011111" => keluaran <= ""; -- -0.58
            when "11111110111011001000011010100011" => keluaran <= ""; -- -0.57
            when "11111110111010010001000000010001" => keluaran <= ""; -- -0.56
            when "11111110111001100001101101001010" => keluaran <= ""; -- -0.55
            when "11111110111000101010010111110010" => keluaran <= ""; -- -0.54
            when "11111110110111110011001010111000" => keluaran <= ""; -- -0.53
            when "11111110110111000000000000010111" => keluaran <= ""; -- -0.52
            when "11111110110110001001010110011100" => keluaran <= ""; -- -0.51
            when "11111110110101010010101010111001" => keluaran <= ""; -- -0.50
            when "11111110110100011100011011110101" => keluaran <= ""; -- -0.49
            when "11111110110011100110011110101011" => keluaran <= ""; -- -0.48
            when "11111110110010110000110111010001" => keluaran <= ""; -- -0.47
            when "11111110110001111111010011001010" => keluaran <= ""; -- -0.46
            when "11111110110001001001101110011011" => keluaran <= ""; -- -0.45
            when "11111110110000010011110011101100" => keluaran <= ""; -- -0.44
            when "11111110101111011101111110100000" => keluaran <= ""; -- -0.43
            when "11111110101110101011110001110001" => keluaran <= ""; -- -0.42
            when "11111110101101110101110110100000" => keluaran <= ""; -- -0.41
            when "11111110101101000000001000011111" => keluaran <= ""; -- -0.40
            when "11111110101100001010011011111110" => keluaran <= ""; -- -0.39
            when "11111110101011010100111111101001" => keluaran <= ""; -- -0.38
            when "11111110101010100011110010011000" => keluaran <= ""; -- -0.37
            when "11111110101001110010101000110111" => keluaran <= ""; -- -0.36
            when "11111110101001000001110101011110" => keluaran <= ""; -- -0.35
            when "11111110101000010001000001101000" => keluaran <= ""; -- -0.34
            when "11111110100111100000000111010101" => keluaran <= ""; -- -0.33
            when "11111110100110110011001100110000" => keluaran <= ""; -- -0.32
            when "11111110100110000010011001100110" => keluaran <= ""; -- -0.31
            when "11111110100101010001110011110001" => keluaran <= ""; -- -0.30
            when "11111110100100100001000111111001" => keluaran <= ""; -- -0.29
            when "11111110100011110000011111100110" => keluaran <= ""; -- -0.28
            when "11111110100011000000000000010000" => keluaran <= ""; -- -0.27
            when "11111110100010010000100110110111" => keluaran <= ""; -- -0.26
            when "11111110100001100001010011000001" => keluaran <= ""; -- -0.25
            when "11111110100000110001101111001000" => keluaran <= ""; -- -0.24
            when "11111110011111111110001000111101" => keluaran <= ""; -- -0.23
            when "11111110011111001110100010010010" => keluaran <= ""; -- -0.22
            when "11111110011110011110111100001011" => keluaran <= ""; -- -0.21
            when "11111110011101101111010010100011" => keluaran <= ""; -- -0.20
            when "11111110011100111111100100110101" => keluaran <= ""; -- -0.19
            when "11111110011011110000000001000011" => keluaran <= ""; -- -0.18
            when "11111110011011000000010110010001" => keluaran <= ""; -- -0.17
            when "11111110011010010000101011010100" => keluaran <= ""; -- -0.16
            when "11111110011001100000111111110110" => keluaran <= ""; -- -0.15
            when "11111110011000110001010100010101" => keluaran <= ""; -- -0.14
            when "11111110010111111101101000010000" => keluaran <= ""; -- -0.13
            when "11111110010111001110000000001010" => keluaran <= ""; -- -0.12
            when "11111110010110011110010011011001" => keluaran <= ""; -- -0.11
            when "11111110010101101110100111001001" => keluaran <= ""; -- -0.10
            when "11111110010100111110111010111101" => keluaran <= ""; -- -0.09
            when "11111110010011101111001110101010" => keluaran <= ""; -- -0.08
            when "11111110010010111110111111011011" => keluaran <= ""; -- -0.07
            when "11111110010010001110110101001000" => keluaran <= ""; -- -0.06
            when "11111110010001011111001011000010" => keluaran <= ""; -- -0.05
            when "11111110010000101111011111110100" => keluaran <= ""; -- -0.04
            when "11111110001111111111110100110001" => keluaran <= ""; -- -0.03
            when "11111110001111001111100011110000" => keluaran <= ""; -- -0.02
            when "11111110001110011111110010100001" => keluaran <= ""; -- -0.01
            when "00000000000000000000000000000000" => keluaran <= ""; --  0.00
            when "00111111011111110000010000011000" => keluaran <= ""; --  0.01
            when "00111111011111100000100000111000" => keluaran <= ""; --  0.02
            when "00111111011111010000110001010000" => keluaran <= ""; --  0.03
            when "00111111011111000001000001101000" => keluaran <= ""; --  0.04
            when "00111111011110110001010010001000" => keluaran <= ""; --  0.05
            when "00111111011110100001100100100000" => keluaran <= ""; --  0.06
            when "00111111011110010001110111100000" => keluaran <= ""; --  0.07
            when "00111111011110000010001001011000" => keluaran <= ""; --  0.08
            when "00111111011101110010011011110000" => keluaran <= ""; --  0.09
            when "00111111011101100010101100101000" => keluaran <= ""; --  0.10
            when "00111111011101010010111101011000" => keluaran <= ""; --  0.11
            when "00111111011101000011001110110000" => keluaran <= ""; --  0.12
            when "00111111011100110011011110001000" => keluaran <= ""; --  0.13
            when "00111111011100100011101111100000" => keluaran <= ""; --  0.14
            when "00111111011011110011111101011000" => keluaran <= ""; --  0.15
            when "00111111011011100011101011110000" => keluaran <= ""; --  0.16
            when "00111111011011010011011010001000" => keluaran <= ""; --  0.17
            when "00111111011011000011001000100000" => keluaran <= ""; --  0.18
            when "00111111011010110010110110111000" => keluaran <= ""; --  0.19
            when "00111111011010100010100101010000" => keluaran <= ""; --  0.20
            when "00111111011010010010010011101000" => keluaran <= ""; --  0.21
            when "00111111011010000010000010000000" => keluaran <= ""; --  0.22
            when "00111111011001110001110000011000" => keluaran <= ""; --  0.23
            when "00111111011001100001100000110000" => keluaran <= ""; --  0.24
            when "00111111011001010001010011001000" => keluaran <= ""; --  0.25
            when "00111111011001000001000100100000" => keluaran <= ""; --  0.26
            when "00111111011000110000110110111000" => keluaran <= ""; --  0.27
            when "00111111011000100000101001010000" => keluaran <= ""; --  0.28
            when "00111111011000010000011111101000" => keluaran <= ""; --  0.29
            when "00111111010111110000010100000000" => keluaran <= ""; --  0.30
            when "00111111010111100000001010011000" => keluaran <= ""; --  0.31
            when "00111111010111010000000000110000" => keluaran <= ""; --  0.32
            when "00111111010111000000010111001000" => keluaran <= ""; --  0.33
            when "00111111010110110000001101111000" => keluaran <= ""; --  0.34
            when "00111111010110100000000011110000" => keluaran <= ""; --  0.35
            when "00111111010110010000011010001000" => keluaran <= ""; --  0.36
            when "00111111010110000000001111111000" => keluaran <= ""; --  0.37
            when "00111111010101110000000101110000" => keluaran <= ""; --  0.38
            when "00111111010101100000011011101000" => keluaran <= ""; --  0.39
            when "00111111010101010000010001110000" => keluaran <= ""; --  0.40
            when "00111111010101000000001011101000" => keluaran <= ""; --  0.41
            when "00111111010100110000000010100000" => keluaran <= ""; --  0.42
            when "00111111010100100000011001011000" => keluaran <= ""; --  0.43
            when "00111111010100010000010000001000" => keluaran <= ""; --  0.44
            when "00111111010011110000000110111000" => keluaran <= ""; --  0.45
            when "00111111010011100000011101110000" => keluaran <= ""; --  0.46
            when "00111111010011010000010100100000" => keluaran <= ""; --  0.47
            when "00111111010011000000001111000000" => keluaran <= ""; --  0.48
            when "00111111010010110000000110010000" => keluaran <= ""; --  0.49
            when "00111111010010100000000001100000" => keluaran <= ""; --  0.50
            when "00111111010010010000011100110000" => keluaran <= ""; --  0.51
            when "00111111010010000000010111011000" => keluaran <= ""; --  0.52
            when "00111111010001110000010010001000" => keluaran <= ""; --  0.53
            when "00111111010001100000001100111000" => keluaran <= ""; --  0.54
            when "00111111010001010000001000001000" => keluaran <= ""; --  0.55
            when "00111111010001000000000011100000" => keluaran <= ""; --  0.56
            when "00111111010000110000000010111000" => keluaran <= ""; --  0.57
            when "00111111010000100000000110010000" => keluaran <= ""; --  0.58
            when "00111111010000010000001001101000" => keluaran <= ""; --  0.59
            when "00111111010000000000001101000000" => keluaran <= ""; --  0.60
            when "00111110111111110000010000011000" => keluaran <= ""; --  0.61
            when "00111110111111100000010000010000" => keluaran <= ""; --  0.62
            when "00111110111111010000010000001000" => keluaran <= ""; --  0.63
            when "00111110111111000000010000000000" => keluaran <= ""; --  0.64
            when "00111110111110110000010000011000" => keluaran <= ""; --  0.65
            when "00111110111110100000010000100000" => keluaran <= ""; --  0.66
            when "00111110111110010000010000101000" => keluaran <= ""; --  0.67
            when "00111110111110000000010000110000" => keluaran <= ""; --  0.68
            when "00111110111101110000010000111000" => keluaran <= ""; --  0.69
            when "00111110111101100000010001000000" => keluaran <= ""; --  0.70
            when "00111110111101010000010001001000" => keluaran <= ""; --  0.71
            when "00111110111101000000010001010000" => keluaran <= ""; --  0.72
            when "00111110111100110000010001011000" => keluaran <= ""; --  0.73
            when "00111110111100100000010001100000" => keluaran <= ""; --  0.74
            when "00111110111100010000010001101000" => keluaran <= ""; --  0.75
            when "00111110111100000000010001110000" => keluaran <= ""; --  0.76
            when "00111110111011110000010001111000" => keluaran <= ""; --  0.77
            when "00111110111011100000010010000000" => keluaran <= ""; --  0.78
            when "00111110111011010000010010001000" => keluaran <= ""; --  0.79
            when "00111110111011000000010010010000" => keluaran <= ""; --  0.80
            when "00111110111010110000010010011000" => keluaran <= ""; --  0.81
            when "00111110111010100000010010100000" => keluaran <= ""; --  0.82
            when "00111110111010010000010010101000" => keluaran <= ""; --  0.83
            when "00111110111010000000010010110000" => keluaran <= ""; --  0.84
            when "00111110111001110000010010111000" => keluaran <= ""; --  0.85
            when "00111110111001100000010011000000" => keluaran <= ""; --  0.86
            when "00111110111001010000010011001000" => keluaran <= ""; --  0.87
            when "00111110111001000000010011010000" => keluaran <= ""; --  0.88
            when "00111110111000110000010011011000" => keluaran <= ""; --  0.89
            when "00111110111000100000010011100000" => keluaran <= ""; --  0.90
            when "00111110111000010000010011101000" => keluaran <= ""; --  0.91
            when "00111110110111110000010100000000" => keluaran <= ""; --  0.92
            when "00111110110111100000010100001000" => keluaran <= ""; --  0.93
            when "00111110110111010000010100010000" => keluaran <= ""; --  0.94
            when "00111110110111000000010100011000" => keluaran <= ""; --  0.95
            when "00111110110110110000010100100000" => keluaran <= ""; --  0.96
            when "00111110110110100000010100101000" => keluaran <= ""; --  0.97
            when "00111110110110010000010100110000" => keluaran <= ""; --  0.98
            when "00111110110110000000010100111000" => keluaran <= ""; --  0.99
            when "00111111100000000000000000000000" => keluaran <= ""; --  1.00
            when others => keluaran <= "0000000000000000";            
        end case;
    end process;
end Behavioral;
